--
-- VHDL Architecture Cursor_test.FSM_test.arch_name
--
-- Created:
--          by - Julie.UNKNOWN (LAPTOP-J400VU4F)
--          at - 12:58:55 10.12.2021
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE arch_name OF FSM_test IS
BEGIN
END ARCHITECTURE arch_name;


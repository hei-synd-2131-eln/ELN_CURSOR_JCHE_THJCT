--
-- VHDL Architecture Cursor_test.Safety_tester.test_safety
--
-- Created:
--          by - Julie.UNKNOWN (LAPTOP-J400VU4F)
--          at - 21:52:41 20.12.2021
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE test_safety OF Safety_tester IS
BEGIN
END ARCHITECTURE test_safety;


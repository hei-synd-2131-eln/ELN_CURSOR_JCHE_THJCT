--
-- VHDL Architecture Cursor_test.Control_DIR_SPEED_tester.test_DIR
--
-- Created:
--          by - Julie.UNKNOWN (LAPTOP-J400VU4F)
--          at - 21:53:55 20.12.2021
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE test_DIR OF Control_DIR_SPEED_tester IS
BEGIN
END ARCHITECTURE test_DIR;

